module test (
    input [2:0] a,
    input [2:0] b,
    output [3:0] c
);
    assign c=a+f+b;
endmodule